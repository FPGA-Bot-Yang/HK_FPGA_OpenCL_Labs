// kernel_system.v

// Generated using ACDS version 17.1.2 304

`timescale 1 ps / 1 ps
module kernel_system (
		input  wire [30:0]  cc_snoop_data,             //          cc_snoop.data
		input  wire         cc_snoop_valid,            //                  .valid
		output wire         cc_snoop_ready,            //                  .ready
		input  wire         cc_snoop_clk_clk,          //      cc_snoop_clk.clk
		input  wire         clock_reset_clk,           //       clock_reset.clk
		input  wire         clock_reset2x_clk,         //     clock_reset2x.clk
		input  wire         clock_reset_reset_reset_n, // clock_reset_reset.reset_n
		output wire         kernel_cra_waitrequest,    //        kernel_cra.waitrequest
		output wire [63:0]  kernel_cra_readdata,       //                  .readdata
		output wire         kernel_cra_readdatavalid,  //                  .readdatavalid
		input  wire [0:0]   kernel_cra_burstcount,     //                  .burstcount
		input  wire [63:0]  kernel_cra_writedata,      //                  .writedata
		input  wire [29:0]  kernel_cra_address,        //                  .address
		input  wire         kernel_cra_write,          //                  .write
		input  wire         kernel_cra_read,           //                  .read
		input  wire [7:0]   kernel_cra_byteenable,     //                  .byteenable
		input  wire         kernel_cra_debugaccess,    //                  .debugaccess
		output wire         kernel_irq_irq,            //        kernel_irq.irq
		input  wire         kernel_mem0_waitrequest,   //       kernel_mem0.waitrequest
		input  wire [511:0] kernel_mem0_readdata,      //                  .readdata
		input  wire         kernel_mem0_readdatavalid, //                  .readdatavalid
		output wire [4:0]   kernel_mem0_burstcount,    //                  .burstcount
		output wire [511:0] kernel_mem0_writedata,     //                  .writedata
		output wire [30:0]  kernel_mem0_address,       //                  .address
		output wire         kernel_mem0_write,         //                  .write
		output wire         kernel_mem0_read,          //                  .read
		output wire [63:0]  kernel_mem0_byteenable,    //                  .byteenable
		output wire         kernel_mem0_debugaccess    //                  .debugaccess
	);

	wire   [63:0] avs_mmm_cra_cra_ring_cra_master_readdata;              // mmm_system:avs_mmm_cra_readdata -> avs_mmm_cra_cra_ring:avm_readdata
	wire          avs_mmm_cra_cra_ring_cra_master_read;                  // avs_mmm_cra_cra_ring:avm_read -> mmm_system:avs_mmm_cra_read
	wire    [3:0] avs_mmm_cra_cra_ring_cra_master_address;               // avs_mmm_cra_cra_ring:avm_addr -> mmm_system:avs_mmm_cra_address
	wire    [7:0] avs_mmm_cra_cra_ring_cra_master_byteenable;            // avs_mmm_cra_cra_ring:avm_byteena -> mmm_system:avs_mmm_cra_byteenable
	wire          avs_mmm_cra_cra_ring_cra_master_readdatavalid;         // mmm_system:avs_mmm_cra_readdatavalid -> avs_mmm_cra_cra_ring:avm_readdatavalid
	wire          avs_mmm_cra_cra_ring_cra_master_write;                 // avs_mmm_cra_cra_ring:avm_write -> mmm_system:avs_mmm_cra_write
	wire   [63:0] avs_mmm_cra_cra_ring_cra_master_writedata;             // avs_mmm_cra_cra_ring:avm_writedata -> mmm_system:avs_mmm_cra_writedata
	wire          clk_1x_out_clk_clk;                                    // clk_1x:out_clk -> [avs_mmm_cra_cra_ring:clk, cra_root:clk, irq_mapper:clk, kernel_cra:clk, kernel_irq:clk, kernel_mem0:clk, mm_interconnect_0:clk_1x_out_clk_clk, mm_interconnect_2:clk_1x_out_clk_clk, mmm_system:clock, reset:clk]
	wire          clk_2x_out_clk_clk;                                    // clk_2x:out_clk -> mmm_system:clock2x
	wire          clk_snoop_out_clk_clk;                                 // clk_snoop:out_clk -> [acl_internal_snoop:in_clk_0_clk, rst_controller:clk]
	wire          avs_mmm_cra_cra_ring_ring_out_datavalid;               // avs_mmm_cra_cra_ring:ro_datavalid -> cra_root:ri_datavalid
	wire          avs_mmm_cra_cra_ring_ring_out_read;                    // avs_mmm_cra_cra_ring:ro_read -> cra_root:ri_read
	wire   [63:0] avs_mmm_cra_cra_ring_ring_out_data;                    // avs_mmm_cra_cra_ring:ro_data -> cra_root:ri_data
	wire    [3:0] avs_mmm_cra_cra_ring_ring_out_addr;                    // avs_mmm_cra_cra_ring:ro_addr -> cra_root:ri_addr
	wire          avs_mmm_cra_cra_ring_ring_out_write;                   // avs_mmm_cra_cra_ring:ro_write -> cra_root:ri_write
	wire    [7:0] avs_mmm_cra_cra_ring_ring_out_byteena;                 // avs_mmm_cra_cra_ring:ro_byteena -> cra_root:ri_byteena
	wire          cra_root_ring_out_datavalid;                           // cra_root:ro_datavalid -> avs_mmm_cra_cra_ring:ri_datavalid
	wire          cra_root_ring_out_read;                                // cra_root:ro_read -> avs_mmm_cra_cra_ring:ri_read
	wire   [63:0] cra_root_ring_out_data;                                // cra_root:ro_data -> avs_mmm_cra_cra_ring:ri_data
	wire    [3:0] cra_root_ring_out_addr;                                // cra_root:ro_addr -> avs_mmm_cra_cra_ring:ri_addr
	wire          cra_root_ring_out_write;                               // cra_root:ro_write -> avs_mmm_cra_cra_ring:ri_write
	wire    [7:0] cra_root_ring_out_byteena;                             // cra_root:ro_byteena -> avs_mmm_cra_cra_ring:ri_byteena
	wire          reset_out_reset_reset;                                 // reset:out_reset_n -> [avs_mmm_cra_cra_ring:rst_n, cra_root:rst_n, irq_mapper:reset, kernel_cra:reset, kernel_irq:reset, kernel_mem0:reset, mm_interconnect_0:mmm_system_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_2:kernel_cra_reset_reset_bridge_in_reset_reset, mmm_system:resetn, rst_controller:reset_in0]
	wire  [511:0] mmm_system_avm_memgmem0_ddr_port_0_0_rw_readdata;      // mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_readdata -> mmm_system:avm_memgmem0_DDR_port_0_0_rw_readdata
	wire          mmm_system_avm_memgmem0_ddr_port_0_0_rw_waitrequest;   // mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_waitrequest -> mmm_system:avm_memgmem0_DDR_port_0_0_rw_waitrequest
	wire   [30:0] mmm_system_avm_memgmem0_ddr_port_0_0_rw_address;       // mmm_system:avm_memgmem0_DDR_port_0_0_rw_address -> mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_address
	wire   [63:0] mmm_system_avm_memgmem0_ddr_port_0_0_rw_byteenable;    // mmm_system:avm_memgmem0_DDR_port_0_0_rw_byteenable -> mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_byteenable
	wire          mmm_system_avm_memgmem0_ddr_port_0_0_rw_read;          // mmm_system:avm_memgmem0_DDR_port_0_0_rw_read -> mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_read
	wire          mmm_system_avm_memgmem0_ddr_port_0_0_rw_readdatavalid; // mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_readdatavalid -> mmm_system:avm_memgmem0_DDR_port_0_0_rw_readdatavalid
	wire          mmm_system_avm_memgmem0_ddr_port_0_0_rw_write;         // mmm_system:avm_memgmem0_DDR_port_0_0_rw_write -> mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_write
	wire  [511:0] mmm_system_avm_memgmem0_ddr_port_0_0_rw_writedata;     // mmm_system:avm_memgmem0_DDR_port_0_0_rw_writedata -> mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_writedata
	wire    [4:0] mmm_system_avm_memgmem0_ddr_port_0_0_rw_burstcount;    // mmm_system:avm_memgmem0_DDR_port_0_0_rw_burstcount -> mm_interconnect_0:mmm_system_avm_memgmem0_DDR_port_0_0_rw_burstcount
	wire  [511:0] mm_interconnect_0_kernel_mem0_s0_readdata;             // kernel_mem0:s0_readdata -> mm_interconnect_0:kernel_mem0_s0_readdata
	wire          mm_interconnect_0_kernel_mem0_s0_waitrequest;          // kernel_mem0:s0_waitrequest -> mm_interconnect_0:kernel_mem0_s0_waitrequest
	wire          mm_interconnect_0_kernel_mem0_s0_debugaccess;          // mm_interconnect_0:kernel_mem0_s0_debugaccess -> kernel_mem0:s0_debugaccess
	wire   [30:0] mm_interconnect_0_kernel_mem0_s0_address;              // mm_interconnect_0:kernel_mem0_s0_address -> kernel_mem0:s0_address
	wire          mm_interconnect_0_kernel_mem0_s0_read;                 // mm_interconnect_0:kernel_mem0_s0_read -> kernel_mem0:s0_read
	wire   [63:0] mm_interconnect_0_kernel_mem0_s0_byteenable;           // mm_interconnect_0:kernel_mem0_s0_byteenable -> kernel_mem0:s0_byteenable
	wire          mm_interconnect_0_kernel_mem0_s0_readdatavalid;        // kernel_mem0:s0_readdatavalid -> mm_interconnect_0:kernel_mem0_s0_readdatavalid
	wire          mm_interconnect_0_kernel_mem0_s0_write;                // mm_interconnect_0:kernel_mem0_s0_write -> kernel_mem0:s0_write
	wire  [511:0] mm_interconnect_0_kernel_mem0_s0_writedata;            // mm_interconnect_0:kernel_mem0_s0_writedata -> kernel_mem0:s0_writedata
	wire    [4:0] mm_interconnect_0_kernel_mem0_s0_burstcount;           // mm_interconnect_0:kernel_mem0_s0_burstcount -> kernel_mem0:s0_burstcount
	wire          kernel_cra_m0_waitrequest;                             // mm_interconnect_2:kernel_cra_m0_waitrequest -> kernel_cra:m0_waitrequest
	wire   [63:0] kernel_cra_m0_readdata;                                // mm_interconnect_2:kernel_cra_m0_readdata -> kernel_cra:m0_readdata
	wire          kernel_cra_m0_debugaccess;                             // kernel_cra:m0_debugaccess -> mm_interconnect_2:kernel_cra_m0_debugaccess
	wire   [29:0] kernel_cra_m0_address;                                 // kernel_cra:m0_address -> mm_interconnect_2:kernel_cra_m0_address
	wire          kernel_cra_m0_read;                                    // kernel_cra:m0_read -> mm_interconnect_2:kernel_cra_m0_read
	wire    [7:0] kernel_cra_m0_byteenable;                              // kernel_cra:m0_byteenable -> mm_interconnect_2:kernel_cra_m0_byteenable
	wire          kernel_cra_m0_readdatavalid;                           // mm_interconnect_2:kernel_cra_m0_readdatavalid -> kernel_cra:m0_readdatavalid
	wire   [63:0] kernel_cra_m0_writedata;                               // kernel_cra:m0_writedata -> mm_interconnect_2:kernel_cra_m0_writedata
	wire          kernel_cra_m0_write;                                   // kernel_cra:m0_write -> mm_interconnect_2:kernel_cra_m0_write
	wire    [0:0] kernel_cra_m0_burstcount;                              // kernel_cra:m0_burstcount -> mm_interconnect_2:kernel_cra_m0_burstcount
	wire   [63:0] mm_interconnect_2_cra_root_cra_slave_readdata;         // cra_root:avs_readdata -> mm_interconnect_2:cra_root_cra_slave_readdata
	wire          mm_interconnect_2_cra_root_cra_slave_waitrequest;      // cra_root:avs_waitrequest -> mm_interconnect_2:cra_root_cra_slave_waitrequest
	wire    [3:0] mm_interconnect_2_cra_root_cra_slave_address;          // mm_interconnect_2:cra_root_cra_slave_address -> cra_root:avs_addr
	wire          mm_interconnect_2_cra_root_cra_slave_read;             // mm_interconnect_2:cra_root_cra_slave_read -> cra_root:avs_read
	wire    [7:0] mm_interconnect_2_cra_root_cra_slave_byteenable;       // mm_interconnect_2:cra_root_cra_slave_byteenable -> cra_root:avs_byteena
	wire          mm_interconnect_2_cra_root_cra_slave_readdatavalid;    // cra_root:avs_readdatavalid -> mm_interconnect_2:cra_root_cra_slave_readdatavalid
	wire          mm_interconnect_2_cra_root_cra_slave_write;            // mm_interconnect_2:cra_root_cra_slave_write -> cra_root:avs_write
	wire   [63:0] mm_interconnect_2_cra_root_cra_slave_writedata;        // mm_interconnect_2:cra_root_cra_slave_writedata -> cra_root:avs_writedata
	wire          irq_mapper_receiver0_irq;                              // mmm_system:kernel_irq -> irq_mapper:receiver0_irq
	wire    [0:0] kernel_irq_receiver_irq_irq;                           // irq_mapper:sender_irq -> kernel_irq:receiver_irq
	wire          rst_controller_reset_out_reset;                        // rst_controller:reset_out -> acl_internal_snoop:in_rst_0_reset

	kernel_system_acl_internal_snoop acl_internal_snoop (
		.in_0_data      (cc_snoop_data),                  //   input,  width = 31,     in_0.data
		.in_0_valid     (cc_snoop_valid),                 //   input,   width = 1,         .valid
		.in_0_ready     (cc_snoop_ready),                 //  output,   width = 1,         .ready
		.in_clk_0_clk   (clk_snoop_out_clk_clk),          //   input,   width = 1, in_clk_0.clk
		.in_rst_0_reset (rst_controller_reset_out_reset), //   input,   width = 1, in_rst_0.reset
		.out_0_data     (),                               //  output,  width = 31,    out_0.data
		.out_0_valid    (),                               //  output,   width = 1,         .valid
		.out_0_ready    ()                                //   input,   width = 1,         .ready
	);

	kernel_system_avs_mmm_cra_cra_ring avs_mmm_cra_cra_ring (
		.clk               (clk_1x_out_clk_clk),                            //   input,   width = 1,      clock.clk
		.avm_read          (avs_mmm_cra_cra_ring_cra_master_read),          //  output,   width = 1, cra_master.read
		.avm_write         (avs_mmm_cra_cra_ring_cra_master_write),         //  output,   width = 1,           .write
		.avm_addr          (avs_mmm_cra_cra_ring_cra_master_address),       //  output,   width = 4,           .address
		.avm_byteena       (avs_mmm_cra_cra_ring_cra_master_byteenable),    //  output,   width = 8,           .byteenable
		.avm_writedata     (avs_mmm_cra_cra_ring_cra_master_writedata),     //  output,  width = 64,           .writedata
		.avm_readdata      (avs_mmm_cra_cra_ring_cra_master_readdata),      //   input,  width = 64,           .readdata
		.avm_readdatavalid (avs_mmm_cra_cra_ring_cra_master_readdatavalid), //   input,   width = 1,           .readdatavalid
		.rst_n             (reset_out_reset_reset),                         //   input,   width = 1,      reset.reset_n
		.ri_read           (cra_root_ring_out_read),                        //   input,   width = 1,    ring_in.read
		.ri_write          (cra_root_ring_out_write),                       //   input,   width = 1,           .write
		.ri_addr           (cra_root_ring_out_addr),                        //   input,   width = 4,           .addr
		.ri_data           (cra_root_ring_out_data),                        //   input,  width = 64,           .data
		.ri_byteena        (cra_root_ring_out_byteena),                     //   input,   width = 8,           .byteena
		.ri_datavalid      (cra_root_ring_out_datavalid),                   //   input,   width = 1,           .datavalid
		.ro_read           (avs_mmm_cra_cra_ring_ring_out_read),            //  output,   width = 1,   ring_out.read
		.ro_write          (avs_mmm_cra_cra_ring_ring_out_write),           //  output,   width = 1,           .write
		.ro_addr           (avs_mmm_cra_cra_ring_ring_out_addr),            //  output,   width = 4,           .addr
		.ro_data           (avs_mmm_cra_cra_ring_ring_out_data),            //  output,  width = 64,           .data
		.ro_byteena        (avs_mmm_cra_cra_ring_ring_out_byteena),         //  output,   width = 8,           .byteena
		.ro_datavalid      (avs_mmm_cra_cra_ring_ring_out_datavalid)        //  output,   width = 1,           .datavalid
	);

	kernel_system_clk_1x clk_1x (
		.in_clk  (clock_reset_clk),    //   input,  width = 1,  in_clk.clk
		.out_clk (clk_1x_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	kernel_system_clk_2x clk_2x (
		.in_clk  (clock_reset2x_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (clk_2x_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	kernel_system_clk_snoop clk_snoop (
		.in_clk  (cc_snoop_clk_clk),      //   input,  width = 1,  in_clk.clk
		.out_clk (clk_snoop_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	kernel_system_cra_root cra_root (
		.clk               (clk_1x_out_clk_clk),                                 //   input,   width = 1,     clock.clk
		.avs_write         (mm_interconnect_2_cra_root_cra_slave_write),         //   input,   width = 1, cra_slave.write
		.avs_addr          (mm_interconnect_2_cra_root_cra_slave_address),       //   input,   width = 4,          .address
		.avs_byteena       (mm_interconnect_2_cra_root_cra_slave_byteenable),    //   input,   width = 8,          .byteenable
		.avs_writedata     (mm_interconnect_2_cra_root_cra_slave_writedata),     //   input,  width = 64,          .writedata
		.avs_readdata      (mm_interconnect_2_cra_root_cra_slave_readdata),      //  output,  width = 64,          .readdata
		.avs_readdatavalid (mm_interconnect_2_cra_root_cra_slave_readdatavalid), //  output,   width = 1,          .readdatavalid
		.avs_waitrequest   (mm_interconnect_2_cra_root_cra_slave_waitrequest),   //  output,   width = 1,          .waitrequest
		.avs_read          (mm_interconnect_2_cra_root_cra_slave_read),          //   input,   width = 1,          .read
		.rst_n             (reset_out_reset_reset),                              //   input,   width = 1,     reset.reset_n
		.ri_write          (avs_mmm_cra_cra_ring_ring_out_write),                //   input,   width = 1,   ring_in.write
		.ri_addr           (avs_mmm_cra_cra_ring_ring_out_addr),                 //   input,   width = 4,          .addr
		.ri_byteena        (avs_mmm_cra_cra_ring_ring_out_byteena),              //   input,   width = 8,          .byteena
		.ri_data           (avs_mmm_cra_cra_ring_ring_out_data),                 //   input,  width = 64,          .data
		.ri_read           (avs_mmm_cra_cra_ring_ring_out_read),                 //   input,   width = 1,          .read
		.ri_datavalid      (avs_mmm_cra_cra_ring_ring_out_datavalid),            //   input,   width = 1,          .datavalid
		.ro_read           (cra_root_ring_out_read),                             //  output,   width = 1,  ring_out.read
		.ro_write          (cra_root_ring_out_write),                            //  output,   width = 1,          .write
		.ro_addr           (cra_root_ring_out_addr),                             //  output,   width = 4,          .addr
		.ro_data           (cra_root_ring_out_data),                             //  output,  width = 64,          .data
		.ro_byteena        (cra_root_ring_out_byteena),                          //  output,   width = 8,          .byteena
		.ro_datavalid      (cra_root_ring_out_datavalid)                         //  output,   width = 1,          .datavalid
	);

	kernel_system_kernel_cra kernel_cra (
		.clk              (clk_1x_out_clk_clk),          //   input,   width = 1,   clk.clk
		.m0_waitrequest   (kernel_cra_m0_waitrequest),   //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (kernel_cra_m0_readdata),      //   input,  width = 64,      .readdata
		.m0_readdatavalid (kernel_cra_m0_readdatavalid), //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (kernel_cra_m0_burstcount),    //  output,   width = 1,      .burstcount
		.m0_writedata     (kernel_cra_m0_writedata),     //  output,  width = 64,      .writedata
		.m0_address       (kernel_cra_m0_address),       //  output,  width = 30,      .address
		.m0_write         (kernel_cra_m0_write),         //  output,   width = 1,      .write
		.m0_read          (kernel_cra_m0_read),          //  output,   width = 1,      .read
		.m0_byteenable    (kernel_cra_m0_byteenable),    //  output,   width = 8,      .byteenable
		.m0_debugaccess   (kernel_cra_m0_debugaccess),   //  output,   width = 1,      .debugaccess
		.reset            (~reset_out_reset_reset),      //   input,   width = 1, reset.reset
		.s0_waitrequest   (kernel_cra_waitrequest),      //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (kernel_cra_readdata),         //  output,  width = 64,      .readdata
		.s0_readdatavalid (kernel_cra_readdatavalid),    //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (kernel_cra_burstcount),       //   input,   width = 1,      .burstcount
		.s0_writedata     (kernel_cra_writedata),        //   input,  width = 64,      .writedata
		.s0_address       (kernel_cra_address),          //   input,  width = 30,      .address
		.s0_write         (kernel_cra_write),            //   input,   width = 1,      .write
		.s0_read          (kernel_cra_read),             //   input,   width = 1,      .read
		.s0_byteenable    (kernel_cra_byteenable),       //   input,   width = 8,      .byteenable
		.s0_debugaccess   (kernel_cra_debugaccess)       //   input,   width = 1,      .debugaccess
	);

	kernel_system_kernel_irq kernel_irq (
		.clk          (clk_1x_out_clk_clk),          //   input,  width = 1,          clk.clk
		.reset        (~reset_out_reset_reset),      //   input,  width = 1,    clk_reset.reset
		.receiver_irq (kernel_irq_receiver_irq_irq), //   input,  width = 1, receiver_irq.irq
		.sender0_irq  (kernel_irq_irq)               //  output,  width = 1,  sender0_irq.irq
	);

	kernel_system_kernel_mem0 kernel_mem0 (
		.clk              (clk_1x_out_clk_clk),                             //   input,    width = 1,   clk.clk
		.m0_waitrequest   (kernel_mem0_waitrequest),                        //   input,    width = 1,    m0.waitrequest
		.m0_readdata      (kernel_mem0_readdata),                           //   input,  width = 512,      .readdata
		.m0_readdatavalid (kernel_mem0_readdatavalid),                      //   input,    width = 1,      .readdatavalid
		.m0_burstcount    (kernel_mem0_burstcount),                         //  output,    width = 5,      .burstcount
		.m0_writedata     (kernel_mem0_writedata),                          //  output,  width = 512,      .writedata
		.m0_address       (kernel_mem0_address),                            //  output,   width = 31,      .address
		.m0_write         (kernel_mem0_write),                              //  output,    width = 1,      .write
		.m0_read          (kernel_mem0_read),                               //  output,    width = 1,      .read
		.m0_byteenable    (kernel_mem0_byteenable),                         //  output,   width = 64,      .byteenable
		.m0_debugaccess   (kernel_mem0_debugaccess),                        //  output,    width = 1,      .debugaccess
		.reset            (~reset_out_reset_reset),                         //   input,    width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_kernel_mem0_s0_waitrequest),   //  output,    width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_kernel_mem0_s0_readdata),      //  output,  width = 512,      .readdata
		.s0_readdatavalid (mm_interconnect_0_kernel_mem0_s0_readdatavalid), //  output,    width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_kernel_mem0_s0_burstcount),    //   input,    width = 5,      .burstcount
		.s0_writedata     (mm_interconnect_0_kernel_mem0_s0_writedata),     //   input,  width = 512,      .writedata
		.s0_address       (mm_interconnect_0_kernel_mem0_s0_address),       //   input,   width = 31,      .address
		.s0_write         (mm_interconnect_0_kernel_mem0_s0_write),         //   input,    width = 1,      .write
		.s0_read          (mm_interconnect_0_kernel_mem0_s0_read),          //   input,    width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_kernel_mem0_s0_byteenable),    //   input,   width = 64,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_kernel_mem0_s0_debugaccess)    //   input,    width = 1,      .debugaccess
	);

	kernel_system_mmm_system mmm_system (
		.avm_mem_gmem0_DDR_port_0_0_rw_address       (mmm_system_avm_memgmem0_ddr_port_0_0_rw_address),       //  output,   width = 31, avm_memgmem0_DDR_port_0_0_rw.address
		.avm_mem_gmem0_DDR_port_0_0_rw_byteenable    (mmm_system_avm_memgmem0_ddr_port_0_0_rw_byteenable),    //  output,   width = 64,                             .byteenable
		.avm_mem_gmem0_DDR_port_0_0_rw_readdatavalid (mmm_system_avm_memgmem0_ddr_port_0_0_rw_readdatavalid), //   input,    width = 1,                             .readdatavalid
		.avm_mem_gmem0_DDR_port_0_0_rw_read          (mmm_system_avm_memgmem0_ddr_port_0_0_rw_read),          //  output,    width = 1,                             .read
		.avm_mem_gmem0_DDR_port_0_0_rw_readdata      (mmm_system_avm_memgmem0_ddr_port_0_0_rw_readdata),      //   input,  width = 512,                             .readdata
		.avm_mem_gmem0_DDR_port_0_0_rw_write         (mmm_system_avm_memgmem0_ddr_port_0_0_rw_write),         //  output,    width = 1,                             .write
		.avm_mem_gmem0_DDR_port_0_0_rw_writedata     (mmm_system_avm_memgmem0_ddr_port_0_0_rw_writedata),     //  output,  width = 512,                             .writedata
		.avm_mem_gmem0_DDR_port_0_0_rw_waitrequest   (mmm_system_avm_memgmem0_ddr_port_0_0_rw_waitrequest),   //   input,    width = 1,                             .waitrequest
		.avm_mem_gmem0_DDR_port_0_0_rw_burstcount    (mmm_system_avm_memgmem0_ddr_port_0_0_rw_burstcount),    //  output,    width = 5,                             .burstcount
		.avs_mmm_cra_read                           (avs_mmm_cra_cra_ring_cra_master_read),                  //   input,    width = 1,                  avs_mmm_cra.read
		.avs_mmm_cra_write                          (avs_mmm_cra_cra_ring_cra_master_write),                 //   input,    width = 1,                             .write
		.avs_mmm_cra_address                        (avs_mmm_cra_cra_ring_cra_master_address),               //   input,    width = 4,                             .address
		.avs_mmm_cra_writedata                      (avs_mmm_cra_cra_ring_cra_master_writedata),             //   input,   width = 64,                             .writedata
		.avs_mmm_cra_byteenable                     (avs_mmm_cra_cra_ring_cra_master_byteenable),            //   input,    width = 8,                             .byteenable
		.avs_mmm_cra_readdata                       (avs_mmm_cra_cra_ring_cra_master_readdata),              //  output,   width = 64,                             .readdata
		.avs_mmm_cra_readdatavalid                  (avs_mmm_cra_cra_ring_cra_master_readdatavalid),         //  output,    width = 1,                             .readdatavalid
		.clock                                      (clk_1x_out_clk_clk),                                    //   input,    width = 1,                  clock_reset.clk
		.clock2x                                    (clk_2x_out_clk_clk),                                    //   input,    width = 1,                clock_reset2x.clk
		.resetn                                     (reset_out_reset_reset),                                 //   input,    width = 1,            clock_reset_reset.reset_n
		.kernel_irq                                 (irq_mapper_receiver0_irq)                               //  output,    width = 1,                   kernel_irq.irq
	);

	kernel_system_reset reset (
		.clk         (clk_1x_out_clk_clk),        //   input,  width = 1,       clk.clk
		.in_reset_n  (clock_reset_reset_reset_n), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (reset_out_reset_reset)      //  output,  width = 1, out_reset.reset_n
	);

	kernel_system_altera_mm_interconnect_171_e6v4f3q mm_interconnect_0 (
		.clk_1x_out_clk_clk                                       (clk_1x_out_clk_clk),                                    //   input,    width = 1,                                     clk_1x_out_clk.clk
		.kernel_mem0_s0_address                                   (mm_interconnect_0_kernel_mem0_s0_address),              //  output,   width = 31,                                     kernel_mem0_s0.address
		.kernel_mem0_s0_write                                     (mm_interconnect_0_kernel_mem0_s0_write),                //  output,    width = 1,                                                   .write
		.kernel_mem0_s0_read                                      (mm_interconnect_0_kernel_mem0_s0_read),                 //  output,    width = 1,                                                   .read
		.kernel_mem0_s0_readdata                                  (mm_interconnect_0_kernel_mem0_s0_readdata),             //   input,  width = 512,                                                   .readdata
		.kernel_mem0_s0_writedata                                 (mm_interconnect_0_kernel_mem0_s0_writedata),            //  output,  width = 512,                                                   .writedata
		.kernel_mem0_s0_burstcount                                (mm_interconnect_0_kernel_mem0_s0_burstcount),           //  output,    width = 5,                                                   .burstcount
		.kernel_mem0_s0_byteenable                                (mm_interconnect_0_kernel_mem0_s0_byteenable),           //  output,   width = 64,                                                   .byteenable
		.kernel_mem0_s0_readdatavalid                             (mm_interconnect_0_kernel_mem0_s0_readdatavalid),        //   input,    width = 1,                                                   .readdatavalid
		.kernel_mem0_s0_waitrequest                               (mm_interconnect_0_kernel_mem0_s0_waitrequest),          //   input,    width = 1,                                                   .waitrequest
		.kernel_mem0_s0_debugaccess                               (mm_interconnect_0_kernel_mem0_s0_debugaccess),          //  output,    width = 1,                                                   .debugaccess
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_address          (mmm_system_avm_memgmem0_ddr_port_0_0_rw_address),       //   input,   width = 31,            mmm_system_avm_memgmem0_DDR_port_0_0_rw.address
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_waitrequest      (mmm_system_avm_memgmem0_ddr_port_0_0_rw_waitrequest),   //  output,    width = 1,                                                   .waitrequest
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_burstcount       (mmm_system_avm_memgmem0_ddr_port_0_0_rw_burstcount),    //   input,    width = 5,                                                   .burstcount
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_byteenable       (mmm_system_avm_memgmem0_ddr_port_0_0_rw_byteenable),    //   input,   width = 64,                                                   .byteenable
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_read             (mmm_system_avm_memgmem0_ddr_port_0_0_rw_read),          //   input,    width = 1,                                                   .read
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_readdata         (mmm_system_avm_memgmem0_ddr_port_0_0_rw_readdata),      //  output,  width = 512,                                                   .readdata
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_readdatavalid    (mmm_system_avm_memgmem0_ddr_port_0_0_rw_readdatavalid), //  output,    width = 1,                                                   .readdatavalid
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_write            (mmm_system_avm_memgmem0_ddr_port_0_0_rw_write),         //   input,    width = 1,                                                   .write
		.mmm_system_avm_memgmem0_DDR_port_0_0_rw_writedata        (mmm_system_avm_memgmem0_ddr_port_0_0_rw_writedata),     //   input,  width = 512,                                                   .writedata
		.mmm_system_clock_reset_reset_reset_bridge_in_reset_reset (~reset_out_reset_reset)                                 //   input,    width = 1, mmm_system_clock_reset_reset_reset_bridge_in_reset.reset
	);

	kernel_system_altera_mm_interconnect_171_w3n7e2q mm_interconnect_2 (
		.clk_1x_out_clk_clk                           (clk_1x_out_clk_clk),                                 //   input,   width = 1,                         clk_1x_out_clk.clk
		.cra_root_cra_slave_address                   (mm_interconnect_2_cra_root_cra_slave_address),       //  output,   width = 4,                     cra_root_cra_slave.address
		.cra_root_cra_slave_write                     (mm_interconnect_2_cra_root_cra_slave_write),         //  output,   width = 1,                                       .write
		.cra_root_cra_slave_read                      (mm_interconnect_2_cra_root_cra_slave_read),          //  output,   width = 1,                                       .read
		.cra_root_cra_slave_readdata                  (mm_interconnect_2_cra_root_cra_slave_readdata),      //   input,  width = 64,                                       .readdata
		.cra_root_cra_slave_writedata                 (mm_interconnect_2_cra_root_cra_slave_writedata),     //  output,  width = 64,                                       .writedata
		.cra_root_cra_slave_byteenable                (mm_interconnect_2_cra_root_cra_slave_byteenable),    //  output,   width = 8,                                       .byteenable
		.cra_root_cra_slave_readdatavalid             (mm_interconnect_2_cra_root_cra_slave_readdatavalid), //   input,   width = 1,                                       .readdatavalid
		.cra_root_cra_slave_waitrequest               (mm_interconnect_2_cra_root_cra_slave_waitrequest),   //   input,   width = 1,                                       .waitrequest
		.kernel_cra_m0_address                        (kernel_cra_m0_address),                              //   input,  width = 30,                          kernel_cra_m0.address
		.kernel_cra_m0_waitrequest                    (kernel_cra_m0_waitrequest),                          //  output,   width = 1,                                       .waitrequest
		.kernel_cra_m0_burstcount                     (kernel_cra_m0_burstcount),                           //   input,   width = 1,                                       .burstcount
		.kernel_cra_m0_byteenable                     (kernel_cra_m0_byteenable),                           //   input,   width = 8,                                       .byteenable
		.kernel_cra_m0_read                           (kernel_cra_m0_read),                                 //   input,   width = 1,                                       .read
		.kernel_cra_m0_readdata                       (kernel_cra_m0_readdata),                             //  output,  width = 64,                                       .readdata
		.kernel_cra_m0_readdatavalid                  (kernel_cra_m0_readdatavalid),                        //  output,   width = 1,                                       .readdatavalid
		.kernel_cra_m0_write                          (kernel_cra_m0_write),                                //   input,   width = 1,                                       .write
		.kernel_cra_m0_writedata                      (kernel_cra_m0_writedata),                            //   input,  width = 64,                                       .writedata
		.kernel_cra_m0_debugaccess                    (kernel_cra_m0_debugaccess),                          //   input,   width = 1,                                       .debugaccess
		.kernel_cra_reset_reset_bridge_in_reset_reset (~reset_out_reset_reset)                              //   input,   width = 1, kernel_cra_reset_reset_bridge_in_reset.reset
	);

	kernel_system_altera_irq_mapper_171_7ezhryi irq_mapper (
		.clk           (clk_1x_out_clk_clk),          //   input,  width = 1,       clk.clk
		.reset         (~reset_out_reset_reset),      //   input,  width = 1, clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),    //   input,  width = 1, receiver0.irq
		.sender_irq    (kernel_irq_receiver_irq_irq)  //  output,  width = 1,    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_out_reset_reset),         //   input,  width = 1, reset_in0.reset
		.clk            (clk_snoop_out_clk_clk),          //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

endmodule
